Miraculous Treasure
aa
